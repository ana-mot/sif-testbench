
package environment_pkg;
    typedef enum {WRITE, READ} direction;
    `include "transaction.svh"
    `include "driver.svh"
    `include "monitor.svh"
endpackage

