package environment_pkg;
    `include "monitor.svh"
endpackage

