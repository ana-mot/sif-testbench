interface reset_if(input logic clk);
  logic rst_b;
endinterface