
package environment_pkg;
    typedef enum {WRITE, READ} direction;
    `include "transaction.svh"
    `include "generator.svh"
    `include "driver.svh"
    `include "monitor.svh"
endpackage

