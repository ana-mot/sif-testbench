
package environment_pkg;
    typedef enum {WRITE, READ} direction;
    `include "transaction.svh"
    `include "generator.svh"
    `include "driver.svh"
    `include "monitor.svh"
    `include "scoreboard.svh"
endpackage

