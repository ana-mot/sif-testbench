class Transaction;
    function new();
        
    endfunction //new()
endclass / Transaction